library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
  port (clk         : in std_logic;
        x           : in unsigned(6 downto 0);
        y           : in unsigned(6 downto 0);
        t_pepe      : in unsigned(3 downto 0);
        data_out    : out std_logic_vector(7 downto 0));
end ram;

architecture Behavioral of ram is
  signal index : unsigned(13 downto 0);

  type ram_t is array (0 to 3599) of std_logic_vector(7 downto 0);
  signal ram : ram_t :=(
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",

x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"72", x"72", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"ba", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba",
x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"72", x"72", x"72", x"72", x"72", x"ba",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"72", x"72", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",

x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba",
x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"ba",
x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"ba",
x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"72", x"72", x"72", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",

x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"ba", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00",
x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"ba", x"72", x"72", x"72", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",

x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"72", x"72", x"72", x"72", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"ba",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba",

x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"ba", x"72", x"72", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"ba", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00",
x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"ba", x"00", x"00", x"00", x"00", x"ba", x"72", x"72", x"ba", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",

x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba",
x"ba", x"72", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"ba",
x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",

x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"ba", x"72", x"72", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",

x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"72", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",

x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba",
x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"72", x"72", x"ba",
x"ba", x"72", x"72", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba",
x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",

x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba",
x"ba", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"ba",
x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",

x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00",
x"ba", x"72", x"72", x"72", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"72", x"ba", x"00", x"00", x"00", x"00", x"00", x"00",
x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"ba", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"


  );
begin
  index <= (to_integer(t_pepe)*300 + y*50 + x);
  process(clk)
  begin
    if rising_edge(clk) then
      data_out <= ram(to_integer(index));
    end if;
  end process;

end Behavioral;
