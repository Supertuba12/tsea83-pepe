library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity scoreMem is
port (
      clk         : in std_logic;
      x           : in unsigned(3 downto 0); -- Range 0 - 15
      y           : in unsigned(3 downto 0); -- Range 0 - 15
      tileIndex   : in unsigned(4 downto 0); -- Range 0 - 17 
      data_out    : out std_logic_vector(7 downto 0));  
end scoreMem;

architecture Behavioral of scoreMem is
  signal index   : unsigned(13 downto 0); -- Change

  type ram_t is array (0 to 4067) of std_logic_vector(7 downto 0);
  signal scoreMem : ram_t :=(
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", -- H
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 

x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", -- I
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 

x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", -- G
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 

x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", -- S
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 

x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", -- C
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 

x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", -- O
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 

x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", -- R
x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 

x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", -- E
x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 

x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", -- 0
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"da", x"da", x"da", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"da", x"da", x"da", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 

x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", -- 1
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 

x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", -- 2
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 

x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", -- 3
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 

x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", -- 4
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 

x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", -- 5
x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 

x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", -- 6
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 

x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", -- 7
x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 

x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", -- 8
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 

x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", -- 9
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"da", x"da", x"da", x"da", x"da", x"da", x"00", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00");

begin  -- scoreMem
  index <= (to_integer(tileIndex*256) + (y*16) + x); -- to_int may not be needed
  data_out <= scoreMem(to_integer(index));

end Behavioral;
 
