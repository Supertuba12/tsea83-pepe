library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ram is
port (
        clk         : in std_logic;
        x           : in integer;
        y           : in integer;
        data_out    : out std_logic_vector(7 downto 0));
end ram;

architecture Behavioral of ram is

    type ram_t is array (0 to 3599) of std_logic_vector(7 downto 0);
    signal ram : ram_t :=(
        x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"70", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 

        x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"70", x"FF", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 

        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"70", 
        x"FF", x"70", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", 
        x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"70", 
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"FF", x"FF", x"FF", 

        x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"70", x"70", x"70", x"FF", 
        x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"70", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"70", x"FF", 
        x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", 
        x"FF", x"FF", x"70", x"70", x"70", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", 

        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", 
        x"70", x"FF", x"70", x"70", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"70", x"FF", x"FF", x"70", x"70", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", 
        x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", 
        x"70", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"70", 
        
        x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"70", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 

        x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"70", x"FF", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 

        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"70", 
        x"FF", x"70", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", 
        x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"70", 
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"FF", x"FF", x"FF", 

        x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"70", x"70", x"70", x"FF", 
        x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"70", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"70", x"FF", 
        x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", 
        x"FF", x"FF", x"70", x"70", x"70", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", 

        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", 
        x"70", x"FF", x"70", x"70", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"70", x"FF", x"FF", x"70", x"70", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", 
        x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", 
        x"70", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"70", 

        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", 
        x"70", x"FF", x"70", x"70", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"70", x"FF", x"FF", x"70", x"70", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", 
        x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", 
        x"70", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"70", 
        
        x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"70", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"70", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"70", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"70", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"70", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"70", x"70", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"

    );
begin
    process(clk)
    begin
        if rising_edge(clk) then
            data_out <= ram(y*50 + x);
        end if;
    end process;    



end Behavioral;
